* Netlist *
C1 2 0 1u
L2 2 3 1u
V3 1 0 1
R4 2 0 100
R5 3 0 100
R6 1 2 100
.end