* Netlist *
C2 2 0 1u
L1 2 3 1u
V2 1 0 1
R2 2 0 100
R3 3 0 100
R1 1 2 100
.end