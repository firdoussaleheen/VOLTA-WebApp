* Translated Netlist *
v V2 1 0
v V1 2 0
q Q1 3 2 0
l L1 1 3
r R1 4 0
c C1 4 0
d D1 3 4
.end