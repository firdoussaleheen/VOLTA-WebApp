*thing*
vAC1 1 0 0 5.00 8000 0 0    
R1 1 0 10ohms
.end
