* Translated Netlist *
v V1 3 0
r R1 4 0
c C1 4 0
d D1 3 4
.end