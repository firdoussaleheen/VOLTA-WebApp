* Netlist *
c C1 2 1 0
l L2 2 1 0
d D1 2 1 0
x X1 3 0 0
q Q1 3 2 0 0 
v V3 1 0 0
r R4 1 2 0
.end
