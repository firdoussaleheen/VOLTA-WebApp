* Translated Netlist *
vV2 1 0
vV1 2 0
qQ1 3 2 0
lL1 1 3
rR1 4 0
cC1 4 0
dD1 3 4
.end