* Translated Netlist *
l L1 V2 Vc
c C1 Vc 0
r R1 Vpulse V2
v V1 Vpulse 0
.end