* Netlist *
C2 2 1 1u
L1 2 1 1u
V2 0 1 1
R1 0 2 100
.end