* Translated Netlist *
v V6 0 5
v V5 6 0
c C2 4 Vout
r R4 4 Vout
r R3 Vout1 4
u U2 Vout 4 0 5 6
v V3 0 3
v V2 1 0
c C1 2 Vout1
r R2 2 Vout1
r R1 Vin 2
v V1 Vin 0
u U1 Vout1 2 0 3 1
.end