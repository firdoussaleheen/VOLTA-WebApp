* Translated Netlist *
v V1 Vac 0
c C1 Vc 0
r R1 Vac Vc
.end